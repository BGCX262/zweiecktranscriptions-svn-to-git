BZh91AY&SYȈ�� ߀Pxg����������`��;�t P.�P�f�I&��h&��5=M<SG�z��@fS���ɢJ�h    h   8i�F#	���12dhh�Q@���Ҁ� 0���db0�`!�M0�!�F��D��&�e=M1MOB2 ���6�*S8DKDh���"FtG0i��Ϋ�����" B��-��~��2	�$N8�!�8�)ä��v.ף!K��|���xy��QN�	��kZx��Q��n�W���c?5cF�hЈ�)IN��Nj�f����:���[��}�ď�I�����u��XpA:ߧh�x�qr�O[D�c�q�Yu`�L5���M�[��2���oQ;1�s&"��:�kgu�Fi�I������g�=/uD3��:�\�ֹq��3j#Y�� m��*���6$�(TӀt[ɲ+��i��%!!!�����A$Y3¶c>���Lgn�%��t��7#�������,@���y��	u�0P�ΈyUd㺿/�����M����
����h�4���߆X6/yY��`�� ���P��F�Kg-Gkf�I���q6G������f�OV�k���u)�q����.W�Wh �����1�䣥qQREW���b�6qB�Q|	�fF�-+�+ZHJ�Ng��;��Vhة�s�T==�7�F�͚�ѳ���Ϊ�u��J��m�H��d�mo2��z��F�#��y�z��<��2�X6�� �q��xS�v�������h��y�9uu3R�E�tu�m_:5���*�����&�>"d.d���f+�o_-��1"An8�B���ޟ3tFc��!V'��x���ZXj���V�fg��ҡ��-��7HE�G@�� f��C��!u�;*�qR�u�;��C����S�i���r���w����7���6�gM��fދ:1\J�u��#�v�5y��1�N8�NJ+����V�c#�9Ery�7s|Z��WW5Xr^mNZ9�A�Q&��ɜ���l8�����d��R����4�	��0�2Qd�) �m��	!!$ܒHD
,���٪��rT���xz"T��FD����B ��	B r�-��+j���@K,�O�.R[}/�ln��.]�HK<X����,�qe-��WH6b�_r�s��#��Ĭ`2������(�\����z#Õ��K���=��]��!Ͽ��"�=�3�[��31����f���kA�:��M� ��$=>A�o�����WS�i#/�<M�א��,ō#�!�l���9Ad�KQڧN�T׳���;Y����uS���ӝR`�8i�M����fA�(7!�jƸ�/�i�	���-�`! �S��>��+��κFl
�Q��J(�n�M�?7%\qL!�M�F{�S^�QGU�78�J��{��Db�i�&n͸>��Vh��g����Y�a�X�<�5'���;�ZP,06""b x���8Q\�N~��Tn �&k ¼�#8E5��+���\(���:�����$p�1)�T�S�����"݊�A�9j�@��:�۫�q�X�I1r٠Έ��Q?T��6^�U�s_ӤfB���9�F�X�"�l�GC%̡�hD
;��c��wl�`�V,��b�8��CQ�y��BI�AӼ�i�X��R�tUx�4T���R��2_�״� )p�Sl��0�3+ɬ5f�C�W!��Q�EЏ<ˏ�D��.<�=��.W�_{A<]w��̹)*~:�=,��&A�7�{�w$S�	��]P